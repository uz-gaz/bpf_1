--------------------------------------------------------------------------------
-- Project Name: A basic processor core for running BPF programs
-- Author:       Fernando Lahoz Bernad
--
-- Description:  Fake instruction RAM for testing. Size: 4096 x 64 bits
--               instructions.
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity Inst_RAM is
    port (
        clk : in std_logic;
        addr : in std_logic_vector (11 downto 0);
        input : in std_logic_vector (63 downto 0);
        write_en : in std_logic;
        read_en : in std_logic;
        output : out std_logic_vector (63 downto 0)
    );
end Inst_RAM;

architecture Behavioral of Inst_RAM is

    type inst_array is array(0 to 4096) of std_logic_vector(63 downto 0);
    signal RAM : inst_array := (
        x"000A0000000001B7",
        x"0000B000000002B7",
        x"00000C00000003B7",
        x"000000D0000004B7",
        x"0000000F000005B7",
        x"0000000000000085",
        x"0000000100000085",
        x"00000010000008B7",
        x"0000000400000837",
        x"0000000200000085",
        x"00000010000008B7",
        x"0000000200000A72",
        x"0000000300000085",
        x"0000000400000085",
        x"0000000500000085",
        x"00010000000001B7",
        x"0000000100000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0002000000000A7A",
        x"000000000000A179",
        x"0000000100000085",
        x"00030000000001B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A279",
        x"0000000100000085",
        x"0000F000000002B7",
        x"00010000000001B7",
        x"0000000200000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0002000000000A7A",
        x"000000000000A179",
        x"0000000200000085",
        x"00030000000001B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A379",
        x"0000000200000085",
        x"000F0000000001B7",
        x"00001000000002B7",
        x"0000000200000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000200000000A7A",
        x"000000000000A279",
        x"0000000200000085",
        x"00003000000002B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A379",
        x"0000000200000085",
        x"0000F000000002B7",
        x"00000F00000003B7",
        x"00010000000001B7",
        x"0000000300000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0002000000000A7A",
        x"000000000000A179",
        x"0000000300000085",
        x"00030000000001B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A479",
        x"0000000300000085",
        x"000F0000000001B7",
        x"00000F00000003B7",
        x"00001000000002B7",
        x"0000000300000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000200000000A7A",
        x"000000000000A279",
        x"0000000300000085",
        x"00003000000002B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A479",
        x"0000000300000085",
        x"000F0000000001B7",
        x"0000F000000002B7",
        x"00000100000003B7",
        x"0000000300000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000020000000A7A",
        x"000000000000A379",
        x"0000000300000085",
        x"00000300000003B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A479",
        x"0000000300000085",
        x"0000F000000002B7",
        x"00000F00000003B7",
        x"000000F0000004B7",
        x"00010000000001B7",
        x"0000000400000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0002000000000A7A",
        x"000000000000A179",
        x"0000000400000085",
        x"00030000000001B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A579",
        x"0000000400000085",
        x"000F0000000001B7",
        x"00000F00000003B7",
        x"000000F0000004B7",
        x"00001000000002B7",
        x"0000000400000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000200000000A7A",
        x"000000000000A279",
        x"0000000400000085",
        x"00003000000002B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A579",
        x"0000000400000085",
        x"000F0000000001B7",
        x"0000F000000002B7",
        x"000000F0000004B7",
        x"00000100000003B7",
        x"0000000400000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000020000000A7A",
        x"000000000000A379",
        x"0000000400000085",
        x"00000300000003B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A579",
        x"0000000400000085",
        x"000F0000000001B7",
        x"0000F000000002B7",
        x"00000F00000003B7",
        x"00000010000004B7",
        x"0000000400000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000002000000A7A",
        x"000000000000A479",
        x"0000000400000085",
        x"00000030000004B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A579",
        x"0000000400000085",
        x"0000F000000002B7",
        x"00000F00000003B7",
        x"000000F0000004B7",
        x"0000000F000005B7",
        x"00010000000001B7",
        x"0000000500000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0002000000000A7A",
        x"000000000000A179",
        x"0000000500000085",
        x"00030000000001B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A679",
        x"0000000500000085",
        x"000F0000000001B7",
        x"00000F00000003B7",
        x"000000F0000004B7",
        x"0000000F000005B7",
        x"00001000000002B7",
        x"0000000500000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000200000000A7A",
        x"000000000000A279",
        x"0000000500000085",
        x"00003000000002B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A679",
        x"0000000500000085",
        x"000F0000000001B7",
        x"0000F000000002B7",
        x"000000F0000004B7",
        x"0000000F000005B7",
        x"00000100000003B7",
        x"0000000500000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000020000000A7A",
        x"000000000000A379",
        x"0000000500000085",
        x"00000300000003B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A679",
        x"0000000500000085",
        x"000F0000000001B7",
        x"0000F000000002B7",
        x"00000F00000003B7",
        x"0000000F000005B7",
        x"00000010000004B7",
        x"0000000500000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000002000000A7A",
        x"000000000000A479",
        x"0000000500000085",
        x"00000030000004B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A679",
        x"0000000500000085",
        x"000F0000000001B7",
        x"0000F000000002B7",
        x"00000F00000003B7",
        x"000000F0000004B7",
        x"00000001000005B7",
        x"0000000500000085",
        x"00000000000008BF",
        x"00000000000009BF",
        x"0000000200000A7A",
        x"000000000000A579",
        x"0000000500000085",
        x"00000003000005B7",
        x"FFFFFFFF00000A7A",
        x"000000000000A679",
        x"0000000500000085",
        x"FFFFFFFF00000085",

        others => x"0000000000000000"
    );

begin

    process (clk)
    begin
        if (clk'event and clk = '1') then
            if (write_en = '1') then
                RAM(conv_integer(addr)) <= input;
            end if;
        end if;
    end process;

    output <= RAM(conv_integer(addr)) when read_en = '1' else (63 downto 0 => '0');

end Behavioral;

