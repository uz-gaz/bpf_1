--------------------------------------------------------------------------------
-- Project Name: A basic processor core for running BPF programs
-- Author:       Fernando Lahoz Bernad
--
-- Description:  Fake instruction RAM for testing. Size: 4096 x 64 bits
--               instructions.
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity Inst_RAM is
    port (
        clk : in std_logic;
        addr : in std_logic_vector (11 downto 0);
        input : in std_logic_vector (63 downto 0);
        write_en : in std_logic;
        read_en : in std_logic;
        output : out std_logic_vector (63 downto 0)
    );
end Inst_RAM;

architecture Behavioral of Inst_RAM is

    type inst_array is array(0 to 4096) of std_logic_vector(63 downto 0);
    signal RAM : inst_array := (
        x"0000000000030005",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"0000000300000006",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"00000018FFFE0815",
        x"00000017000009B7",
        x"000000000003981D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"00000017FFFE0855",
        x"00000018000009B7",
        x"000000000003985D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"00000017FFFE0825",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000FFFB982D",
        x"00000010000008B7",
        x"00000007000009B7",
        x"000000000003982D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"0000001700030835",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000FFFD983D",
        x"00000010000008B7",
        x"00000007000009B7",
        x"000000000003983D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"00000017FFFE0865",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000FFFB986D",
        x"00000010000008B7",
        x"00000007000009B7",
        x"000000000003986D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFE9000008B7",
        x"FFFFFFEF000009B7",
        x"00000000FFFD986D",
        x"FFFFFFD6000008B7",
        x"FFFFFFCC00030865",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"0000001700030875",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000FFFD987D",
        x"00000010000008B7",
        x"00000007000009B7",
        x"000000000003987D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFE9000008B7",
        x"FFFFFFEF000009B7",
        x"00000000FFFD987D",
        x"FFFFFFD6000008B7",
        x"FFFFFFCC00030875",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000017000008B7",
        x"00000017FFFE08A5",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000000398AD",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000010000008B7",
        x"00000007000009B7",
        x"00000000FFFD98AD",
        x"00000017000008B7",
        x"00000017000308B5",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000000398BD",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000010000008B7",
        x"00000007000009B7",
        x"00000000FFFD98BD",
        x"00000017000008B7",
        x"00000017000608C5",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000000398CD",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000010000008B7",
        x"00000007000009B7",
        x"00000000FFFD98CD",
        x"FFFFFFE9000008B7",
        x"FFFFFFEF000009B7",
        x"00000000000398CD",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFD6000008B7",
        x"FFFFFFCCFFFE08C5",
        x"00000017000008B7",
        x"00000017000308D5",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"0000000E000008B7",
        x"0000000F000009B7",
        x"00000000000398DD",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000010000008B7",
        x"00000007000009B7",
        x"00000000FFFD98DD",
        x"FFFFFFE9000008B7",
        x"FFFFFFEF000009B7",
        x"00000000000398CD",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFD6000008B7",
        x"FFFFFFCCFFFE08C5",
        x"0000000000040005",
        x"0000000000000095",
        x"FFFFFFFE000000B7",
        x"FFFFFFFE000001B7",
        x"FFFFFFFE000002B7",
        x"00000017000008B7",
        x"0000000100030845",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"00000008000008B7",
        x"00000004000009B7",
        x"00000000FFFD984D",
        x"FFFFFFFF000008B7",
        x"0000004B000009B7",
        x"000000000003984D",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFE9000008B4",
        x"FFFFFFEF000009B4",
        x"00000000FFFD986E",
        x"FFFFFFD6000008B4",
        x"FFFFFFCC00030866",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFE9000008B4",
        x"FFFFFFEF000009B4",
        x"00000000FFFD987D",
        x"FFFFFFD6000008B4",
        x"FFFFFFCC00030876",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFE9000008B4",
        x"FFFFFFEF000009B4",
        x"00000000000398CE",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFD6000008B4",
        x"FFFFFFCCFFFE08C6",
        x"FFFFFFE9000008B4",
        x"FFFFFFEF000009B4",
        x"00000000000398CE",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",
        x"FFFFFFD6000008B4",
        x"FFFFFFCCFFFE08C6",
        x"000000000001001D",
        x"000000000003111D",
        x"000000000001221D",
        x"000000000001331D",
        x"00000000FFC90005",
        x"FFFFFFFF000000B7",
        x"FFFFFFFF000001B7",
        x"FFFFFFFF000002B7",

        others => x"0000000000000000"
    );

begin

    process (clk)
    begin
        if (clk'event and clk = '1') then
            if (write_en = '1') then
                RAM(conv_integer(addr)) <= input;
            end if;
        end if;
    end process;

    output <= RAM(conv_integer(addr)) when read_en = '1' else (63 downto 0 => '0');

end Behavioral;

