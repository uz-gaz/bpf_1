--------------------------------------------------------------------------------
-- Project Name: A basic processor core for running BPF programs
-- Author:       Fernando Lahoz Bernad
--
-- Description:  Fake instruction RAM for testing. Size: 4096 x 64 bits
--               instructions.
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity Inst_RAM is
    port (
        clk : in std_logic;
        addr : in std_logic_vector (11 downto 0);
        input : in std_logic_vector (63 downto 0);
        write_en : in std_logic;
        read_en : in std_logic;
        output : out std_logic_vector (63 downto 0)
    );
end Inst_RAM;

architecture Behavioral of Inst_RAM is

    type inst_array is array(0 to 4096) of std_logic_vector(63 downto 0);
    signal RAM : inst_array := (
        x"0000004000000607",
        x"000000000000460F",
        x"0000004000000617",
        x"000000000000461F",
        x"0000004000000627",
        x"000000000000462F",
        x"0000004000000637",
        x"000000000000463F",
        x"0000004000010637",
        x"000000000001463F",
        x"0000004000000647",
        x"000000000000464F",
        x"0000004000000657",
        x"000000000000465F",
        x"0000004000000667",
        x"000000000000466F",
        x"0000004000000677",
        x"000000000000467F",
        x"0000000000000687",
        x"0000004000000697",
        x"000000000000469F",
        x"0000004000010697",
        x"000000000001469F",
        x"00000040000006A7",
        x"00000000000046AF",
        x"00000040000006B7",
        x"00000000000046BF",
        x"00000040000806B7",
        x"00000000000846BF",
        x"00000040001006B7",
        x"00000000001046BF",
        x"00000040002006B7",
        x"00000000002046BF",
        x"00000040000006C7",
        x"00000000000046CF",
        x"0000002000000304",
        x"000000000000230C",
        x"0000002000000314",
        x"000000000000231C",
        x"0000002000000324",
        x"000000000000232C",
        x"0000002000000334",
        x"000000000000233C",
        x"0000002000010334",
        x"000000000001233C",
        x"0000002000000344",
        x"000000000000234C",
        x"0000002000000354",
        x"000000000000235C",
        x"0000002000000364",
        x"000000000000236C",
        x"0000002000000374",
        x"000000000000237C",
        x"0000000000000384",
        x"0000002000000394",
        x"000000000000239C",
        x"0000002000010394",
        x"000000000001239C",
        x"00000020000003A4",
        x"00000000000023AC",
        x"00000020000003B4",
        x"00000000000023BC",
        x"00000020000803B4",
        x"00000000000823BC",
        x"00000020001003B4",
        x"00000000001023BC",
        x"00000020000003C4",
        x"00000000000023CC",
        x"00000010000007D4",
        x"00000020000007D4",
        x"00000040000007D4",
        x"00000010000007DC",
        x"00000020000007DC",
        x"00000040000007DC",
        x"00000010000007D7",
        x"00000020000007D7",
        x"00000040000007D7",
        x"00000000003651C3",
        x"00000000003651DB",
        x"00000050003651C3",
        x"00000050003651DB",
        x"00000040003651C3",
        x"00000040003651DB",
        x"000000A0003651C3",
        x"000000A0003651DB",
        x"00000001003651C3",
        x"00000001003651DB",
        x"00000051003651C3",
        x"00000051003651DB",
        x"00000041003651C3",
        x"00000041003651DB",
        x"000000A1003651C3",
        x"000000A1003651DB",
        x"000000E1003651C3",
        x"000000E1003651DB",
        x"000000F1003651C3",
        x"000000F1003651DB",
        x"FFFFFFF600000718",
        x"FFFFFFFF00000000",
        x"0000000000659771",
        x"0000000000659769",
        x"0000000000659761",
        x"0000000000659779",
        x"0000000000659789",
        x"0000000000659791",
        x"0000000000659781",
        x"0000005000650772",
        x"000000500065076A",
        x"0000005000650762",
        x"000000500065077A",
        x"0000000000659773",
        x"000000000065976B",
        x"0000000000659763",
        x"000000000065977B",
        x"0000000000000005",
        x"0000000C00000115",
        x"000000000000A11D",
        x"0000000C00000125",
        x"000000000000A12D",
        x"0000000C00000135",
        x"000000000000A13D",
        x"0000000C000001A5",
        x"000000000000A1AD",
        x"0000000C000001B5",
        x"000000000000A1BD",
        x"0000000C00000145",
        x"000000000000A14D",
        x"0000000C00000155",
        x"000000000000A15D",
        x"0000000C00000165",
        x"000000000000A16D",
        x"0000000C00000175",
        x"000000000000A17D",
        x"0000000C000001C5",
        x"000000000000A1CD",
        x"0000000C000001D5",
        x"000000000000A1DD",
        x"0000000C00000085",
        x"0000000000000006",
        x"0000000C00000116",
        x"000000000000A11E",
        x"0000000C00000126",
        x"000000000000A12E",
        x"0000000C00000136",
        x"000000000000A13E",
        x"0000000C000001A6",
        x"000000000000A1AE",
        x"0000000C000001B6",
        x"000000000000A1BE",
        x"0000000C00000146",
        x"000000000000A14E",
        x"0000000C00000156",
        x"000000000000A15E",
        x"0000000C00000166",
        x"000000000000A16E",
        x"0000000C00000176",
        x"000000000000A17E",
        x"0000000C000001C6",
        x"000000000000A1CE",
        x"0000000C000001D6",
        x"000000000000A1DE",
        x"0000000000000095",

        others => x"0000000000000000"
    );

begin

    process (clk)
    begin
        if (clk'event and clk = '1') then
            if (write_en = '1') then
                RAM(conv_integer(addr)) <= input;
            end if;
        end if;
    end process;

    output <= RAM(conv_integer(addr)) when read_en = '1' else (63 downto 0 => '0');

end Behavioral;